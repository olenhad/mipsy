----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    10:52:17 10/23/2013 
-- Design Name: 
-- Module Name:    funct_to_alu - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity funct_to_alu is
	Port ( funct : in  STD_LOGIC_VECTOR(5 downto 0);
			 alu_ctrl : out std_logic_vector(5 downto 0));
end funct_to_alu;

architecture Behavioral of funct_to_alu is

begin

alu_ctrl <= 

end Behavioral;

