x"01", x"10", x"01", x"3c", x"00", x"00", x"29", x"8c", x"01", x"10", x"01", x"3c", x"04", x"00", x"2a", x"8c", 
x"20", x"58", x"49", x"01", x"01", x"10", x"01", x"3c", x"3c", x"00", x"2b", x"ac", x"07", x"00", x"10", x"08", 
