x"01", x"10", x"01", x"3c", x"00", x"00", x"29", x"8c", x"01", x"10", x"01", x"3c", x"04", x"00", x"2a", x"8c", 
x"20", x"58", x"49", x"01", x"22", x"78", x"69", x"01", x"01", x"10", x"01", x"3c", x"08", x"00", x"29", x"8c", 
x"01", x"00", x"e9", x"11", x"09", x"00", x"10", x"08", x"01", x"10", x"01", x"3c", x"3c", x"00", x"2f", x"ac", 
x"09", x"00", x"10", x"08", 